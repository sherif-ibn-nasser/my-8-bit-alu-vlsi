magic
tech scmos
timestamp 1734629465
<< ndiffusion >>
rect 65 19 66 23
rect 503 19 504 23
<< metal1 >>
rect 0 65 52 69
rect 74 65 490 69
rect 512 65 568 69
rect 590 65 615 69
rect 66 30 70 37
rect 481 29 497 33
rect 504 30 508 37
rect 66 23 70 26
rect 566 29 575 33
rect 619 32 622 36
rect 504 23 508 26
rect 0 5 52 9
rect 65 5 71 9
rect 74 5 490 9
rect 512 5 568 9
rect 590 5 615 9
<< metal2 >>
rect -7 65 -4 69
rect 66 30 70 32
rect 461 29 477 33
rect 504 30 508 32
rect 551 29 562 33
rect 611 32 615 36
rect 582 30 586 32
rect 623 24 629 28
<< metal3 >>
rect -12 69 -6 74
rect -12 65 -11 69
rect -7 65 -6 69
rect -12 5 -6 65
rect 22 5 28 74
rect 65 36 71 37
rect 65 32 66 36
rect 70 32 71 36
rect 65 5 71 32
rect 105 5 111 74
rect 456 33 462 74
rect 456 29 457 33
rect 461 29 462 33
rect 456 5 462 29
rect 503 36 509 37
rect 503 32 504 36
rect 508 32 509 36
rect 503 5 509 32
rect 546 33 552 74
rect 546 29 547 33
rect 551 29 552 33
rect 546 5 552 29
rect 581 36 587 37
rect 581 32 582 36
rect 586 32 587 36
rect 581 5 587 32
rect 606 36 612 74
rect 606 32 607 36
rect 611 32 612 36
rect 606 5 612 32
rect 618 28 624 29
rect 618 24 619 28
rect 623 24 624 28
rect 618 5 624 24
<< polycontact >>
rect 497 29 501 33
rect 575 29 579 33
rect 622 32 626 36
<< ndcontact >>
rect 66 19 70 23
rect 504 19 508 23
<< m2contact >>
rect -4 65 0 69
rect 66 26 70 30
rect 477 29 481 33
rect 504 26 508 30
rect 562 29 566 33
rect 615 32 619 36
rect 582 26 586 30
rect 629 24 633 28
<< m3contact >>
rect -11 65 -7 69
rect 66 32 70 36
rect 457 29 461 33
rect 504 32 508 36
rect 547 29 551 33
rect 582 32 586 36
rect 607 32 611 36
rect 619 24 623 28
use inv  inv_0
timestamp 1734626176
transform 1 0 52 0 1 19
box 0 -14 22 50
use inv  inv_1
timestamp 1734626176
transform 1 0 615 0 1 19
box 0 -14 22 50
use inv  inv_2
timestamp 1734626176
transform 1 0 490 0 1 19
box 0 -14 22 50
use inv  inv_3
timestamp 1734626176
transform 1 0 568 0 1 19
box 0 -14 22 50
<< labels >>
flabel metal3 -10 69 -6 74 0 FreeMono 40 0 0 0 VDD
port 1 nsew
flabel metal3 22 69 28 74 0 FreeMono 40 0 0 0 InvB
port 3 nsew
flabel metal3 105 69 111 74 0 FreeMono 40 0 0 0 GND
port 5 nsew
flabel metal3 456 69 462 74 0 FreeMono 40 0 0 0 OP0
port 7 nsew
flabel metal3 546 69 552 74 0 FreeMono 40 0 0 0 OP1
port 9 nsew
flabel metal3 606 69 612 74 0 FreeMono 40 0 0 0 InvOut
port 11 nsew
<< end >>
