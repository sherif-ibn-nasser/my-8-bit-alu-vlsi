magic
tech scmos
timestamp 1734627670
<< nwell >>
rect 0 20 32 40
<< polysilicon >>
rect 9 36 13 42
rect 19 36 23 42
rect 9 4 13 24
rect 19 4 23 24
rect 9 -6 13 0
rect 19 -6 23 0
<< ndiffusion >>
rect 8 0 9 4
rect 13 0 14 4
rect 18 0 19 4
rect 23 0 24 4
<< pdiffusion >>
rect 8 24 9 36
rect 13 24 19 36
rect 23 24 24 36
<< metal1 >>
rect 0 46 32 50
rect 4 36 8 46
rect 24 16 28 24
rect 14 12 28 16
rect 14 4 18 12
rect 4 -10 8 0
rect 24 -10 28 0
rect 0 -14 32 -10
<< ntransistor >>
rect 9 0 13 4
rect 19 0 23 4
<< ptransistor >>
rect 9 24 13 36
rect 19 24 23 36
<< ndcontact >>
rect 4 0 8 4
rect 14 0 18 4
rect 24 0 28 4
<< pdcontact >>
rect 4 24 8 36
rect 24 24 28 36
<< labels >>
flabel metal1 0 46 32 50 0 FreeMono 40 0 0 0 VDD
port 1 nsew
flabel metal1 0 -14 32 -10 0 FreeMono 40 0 0 0 GND
port 3 nsew
flabel polysilicon 9 -6 13 -2 0 FreeMono 40 0 0 0 X
port 5 nsew
flabel polysilicon 19 -6 23 -2 0 FreeMono 40 0 0 0 Y
port 6 nsew
<< end >>
